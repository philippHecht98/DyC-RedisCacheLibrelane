package cache_cfg_pkg;

    localparam int unsigned NUM_ENTRIES = 16;
    localparam int unsigned KEY_WIDTH   = 32;
    localparam int unsigned VALUE_WIDTH = 64;

endpackage